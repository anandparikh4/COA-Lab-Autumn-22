`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:08:15 09/13/2022 
// Design Name: 
// Module Name:    Q2_Grp_81 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Q2_Grp_81(input [3:0] counter,output [3:0] sum, output carry);
wire c0,c1,c2;


endmodule
